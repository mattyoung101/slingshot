module mod (
    input logic foo1,
    output logic foo2
);
    assign foo1 = foo2;
endmodule
